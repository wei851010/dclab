// lab2.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module lab2 (
		input  wire  clk_clk,                        //                        clk.clk
		input  wire  reset_reset_n,                  //                      reset.reset_n
		input  wire  uart_0_external_connection_RXD, // uart_0_external_connection.RXD
		output wire  uart_0_external_connection_TXD  //                           .TXD
	);

	wire         altpll_0_c0_clk;                                         // altpll_0:c0 -> [Rsa256Wrapper_0:avm_clk, mm_interconnect_0:altpll_0_c0_clk, rs232_0:clk, rst_controller:clk]
	wire  [31:0] rsa256wrapper_0_avalon_master_0_readdata;                // mm_interconnect_0:Rsa256Wrapper_0_avalon_master_0_readdata -> Rsa256Wrapper_0:avm_readdata
	wire         rsa256wrapper_0_avalon_master_0_waitrequest;             // mm_interconnect_0:Rsa256Wrapper_0_avalon_master_0_waitrequest -> Rsa256Wrapper_0:avm_waitrequest
	wire   [4:0] rsa256wrapper_0_avalon_master_0_address;                 // Rsa256Wrapper_0:avm_address -> mm_interconnect_0:Rsa256Wrapper_0_avalon_master_0_address
	wire         rsa256wrapper_0_avalon_master_0_read;                    // Rsa256Wrapper_0:avm_read -> mm_interconnect_0:Rsa256Wrapper_0_avalon_master_0_read
	wire         rsa256wrapper_0_avalon_master_0_write;                   // Rsa256Wrapper_0:avm_write -> mm_interconnect_0:Rsa256Wrapper_0_avalon_master_0_write
	wire  [31:0] rsa256wrapper_0_avalon_master_0_writedata;               // Rsa256Wrapper_0:avm_writedata -> mm_interconnect_0:Rsa256Wrapper_0_avalon_master_0_writedata
	wire         mm_interconnect_0_rs232_0_avalon_rs232_slave_chipselect; // mm_interconnect_0:rs232_0_avalon_rs232_slave_chipselect -> rs232_0:chipselect
	wire  [31:0] mm_interconnect_0_rs232_0_avalon_rs232_slave_readdata;   // rs232_0:readdata -> mm_interconnect_0:rs232_0_avalon_rs232_slave_readdata
	wire   [0:0] mm_interconnect_0_rs232_0_avalon_rs232_slave_address;    // mm_interconnect_0:rs232_0_avalon_rs232_slave_address -> rs232_0:address
	wire         mm_interconnect_0_rs232_0_avalon_rs232_slave_read;       // mm_interconnect_0:rs232_0_avalon_rs232_slave_read -> rs232_0:read
	wire   [3:0] mm_interconnect_0_rs232_0_avalon_rs232_slave_byteenable; // mm_interconnect_0:rs232_0_avalon_rs232_slave_byteenable -> rs232_0:byteenable
	wire         mm_interconnect_0_rs232_0_avalon_rs232_slave_write;      // mm_interconnect_0:rs232_0_avalon_rs232_slave_write -> rs232_0:write
	wire  [31:0] mm_interconnect_0_rs232_0_avalon_rs232_slave_writedata;  // mm_interconnect_0:rs232_0_avalon_rs232_slave_writedata -> rs232_0:writedata
	wire         rst_controller_reset_out_reset;                          // rst_controller:reset_out -> [Rsa256Wrapper_0:avm_rst, mm_interconnect_0:Rsa256Wrapper_0_reset_sink_reset_bridge_in_reset_reset, rs232_0:reset]
	wire         rst_controller_001_reset_out_reset;                      // rst_controller_001:reset_out -> altpll_0:reset

	Rsa256Wrapper rsa256wrapper_0 (
		.avm_address     (rsa256wrapper_0_avalon_master_0_address),     // avalon_master_0.address
		.avm_read        (rsa256wrapper_0_avalon_master_0_read),        //                .read
		.avm_readdata    (rsa256wrapper_0_avalon_master_0_readdata),    //                .readdata
		.avm_write       (rsa256wrapper_0_avalon_master_0_write),       //                .write
		.avm_writedata   (rsa256wrapper_0_avalon_master_0_writedata),   //                .writedata
		.avm_waitrequest (rsa256wrapper_0_avalon_master_0_waitrequest), //                .waitrequest
		.avm_clk         (altpll_0_c0_clk),                             //      clock_sink.clk
		.avm_rst         (rst_controller_reset_out_reset)               //      reset_sink.reset
	);

	lab2_altpll_0 altpll_0 (
		.clk       (clk_clk),                            //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset), // inclk_interface_reset.reset
		.read      (),                                   //             pll_slave.read
		.write     (),                                   //                      .write
		.address   (),                                   //                      .address
		.readdata  (),                                   //                      .readdata
		.writedata (),                                   //                      .writedata
		.c0        (altpll_0_c0_clk),                    //                    c0.clk
		.areset    (),                                   //        areset_conduit.export
		.locked    (),                                   //        locked_conduit.export
		.phasedone ()                                    //     phasedone_conduit.export
	);

	lab2_rs232_0 rs232_0 (
		.clk        (altpll_0_c0_clk),                                         //                clk.clk
		.reset      (rst_controller_reset_out_reset),                          //              reset.reset
		.address    (mm_interconnect_0_rs232_0_avalon_rs232_slave_address),    // avalon_rs232_slave.address
		.chipselect (mm_interconnect_0_rs232_0_avalon_rs232_slave_chipselect), //                   .chipselect
		.byteenable (mm_interconnect_0_rs232_0_avalon_rs232_slave_byteenable), //                   .byteenable
		.read       (mm_interconnect_0_rs232_0_avalon_rs232_slave_read),       //                   .read
		.write      (mm_interconnect_0_rs232_0_avalon_rs232_slave_write),      //                   .write
		.writedata  (mm_interconnect_0_rs232_0_avalon_rs232_slave_writedata),  //                   .writedata
		.readdata   (mm_interconnect_0_rs232_0_avalon_rs232_slave_readdata),   //                   .readdata
		.irq        (),                                                        //          interrupt.irq
		.UART_RXD   (uart_0_external_connection_RXD),                          // external_interface.export
		.UART_TXD   (uart_0_external_connection_TXD)                           //                   .export
	);

	lab2_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                        (altpll_0_c0_clk),                                         //                                      altpll_0_c0.clk
		.Rsa256Wrapper_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                          // Rsa256Wrapper_0_reset_sink_reset_bridge_in_reset.reset
		.Rsa256Wrapper_0_avalon_master_0_address                (rsa256wrapper_0_avalon_master_0_address),                 //                  Rsa256Wrapper_0_avalon_master_0.address
		.Rsa256Wrapper_0_avalon_master_0_waitrequest            (rsa256wrapper_0_avalon_master_0_waitrequest),             //                                                 .waitrequest
		.Rsa256Wrapper_0_avalon_master_0_read                   (rsa256wrapper_0_avalon_master_0_read),                    //                                                 .read
		.Rsa256Wrapper_0_avalon_master_0_readdata               (rsa256wrapper_0_avalon_master_0_readdata),                //                                                 .readdata
		.Rsa256Wrapper_0_avalon_master_0_write                  (rsa256wrapper_0_avalon_master_0_write),                   //                                                 .write
		.Rsa256Wrapper_0_avalon_master_0_writedata              (rsa256wrapper_0_avalon_master_0_writedata),               //                                                 .writedata
		.rs232_0_avalon_rs232_slave_address                     (mm_interconnect_0_rs232_0_avalon_rs232_slave_address),    //                       rs232_0_avalon_rs232_slave.address
		.rs232_0_avalon_rs232_slave_write                       (mm_interconnect_0_rs232_0_avalon_rs232_slave_write),      //                                                 .write
		.rs232_0_avalon_rs232_slave_read                        (mm_interconnect_0_rs232_0_avalon_rs232_slave_read),       //                                                 .read
		.rs232_0_avalon_rs232_slave_readdata                    (mm_interconnect_0_rs232_0_avalon_rs232_slave_readdata),   //                                                 .readdata
		.rs232_0_avalon_rs232_slave_writedata                   (mm_interconnect_0_rs232_0_avalon_rs232_slave_writedata),  //                                                 .writedata
		.rs232_0_avalon_rs232_slave_byteenable                  (mm_interconnect_0_rs232_0_avalon_rs232_slave_byteenable), //                                                 .byteenable
		.rs232_0_avalon_rs232_slave_chipselect                  (mm_interconnect_0_rs232_0_avalon_rs232_slave_chipselect)  //                                                 .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (altpll_0_c0_clk),                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
