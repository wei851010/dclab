
module lab2 (
	clk_clk,
	reset_reset_n,
	uart_0_external_connection_RXD,
	uart_0_external_connection_TXD);	

	input		clk_clk;
	input		reset_reset_n;
	input		uart_0_external_connection_RXD;
	output		uart_0_external_connection_TXD;
endmodule
